4,8,QR���`��,Q,113,,0,0 01 00 0,113,6661736B646C666A61736A64666C6B616A7364666C6B6A61736C646A6B663B6C6173646A666C3B61736B6A64663B6C61736A6B64666C3B61736A64663B6C61736B6A64676B6864736A6B66676B6A73646866676B6A73646B666A67686B73646A66676B6C6A73646C6B66676A6C73646667,,,,,,
