4,8,QR���`��,Q,43,,0,0 01 00 0,43,687474703A2F2F77656978696E2E71712E636F6D2F722F4E485561416A33455F47434872586C683979416D,,,,,,
