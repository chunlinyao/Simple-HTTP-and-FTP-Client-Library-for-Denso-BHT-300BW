4,8,QR���`��,Q,20,,0,0 01 00 0,20,315053323543333330484353342D412B43333235,,,,,,
4,8,QR���`��,Q,37,,0,0 01 00 0,37,51523153364B31303030304843352A30303230302A353031365431392A35302A36302A2A2A,,,,,,
4,8,QR���`��,Q,37,,0,0 01 00 0,37,51523153313053453130304653352A30303230302A363231355433332A35302A36302A2A2A,,,,,,
4,4,CODE39,M,8,1T506T8Z,0,,8,315435303654385A,,,,,,
4,8,QR���`��,Q,4,,0,0 01 00 0,4,51333435,,,,,,
4,8,QR���`��,Q,5,,0,0 01 00 0,5,433A4F5054,,,,,,
4,8,QR���`��,Q,6,,0,0 01 00 0,6,504C543A3333,,,,,,
4,8,QR���`��,Q,5,,0,0 01 00 0,5,433A334445,,,,,,
4,8,QR���`��,Q,6,,0,0 01 00 0,6,504C543A3230,,,,,,
4,8,QR���`��,Q,5,,0,0 01 00 0,5,433A414944,,,,,,
4,8,QR���`��,Q,11,,0,0 01 00 0,11,31506E6F74657869737473,,,,,,
